VS1  VDD 0 DC 5
VS2  q1b 0 PULSE(0 5 0 0 0 5m 20m)
VS3  q2b 0 PULSE(0 5 10m 0 0 5m 20m)


R1  q1c vdd 1k
Q1  q1c q1b 0 QNPN
R2  q1b q2c 10k

R3  q2c vdd 1k
Q2  q2c q2b 0 QNPN
R4  q2b q1c 10k

*bc547b
.MODEL QNPN  NPN (BF=530 NE=1.3 ISE=9.72F IKF=80M IS=20F VAF=50V
+      BR=10 NC=2 ISC=47P IKR=12M VAR=10
+      RB=280 RE=1 RC=40 TR=.3U
+      CJE=12P VJE=.48 MJE=0.5 CJC=6P VJC=.7 MJC=.33 TF=.5N)

.TRAN .1m 100m 

.end