VS1  VDD 0 DC 5
VS2  nor1b 0 DC 0
*PULSE(0 5 1n 0 0 5m 20m)
VS3  nor2b 0 DC 0
*PULSE(0 5 10.001m 0 0 5m 20m)
*init sr latch
VS4  nor1q 0 PULSE(0 5 0 0 0 1n 0)

*nor 1
Q1  nor1q nor1a 0 QNPN
Q2  nor1q nor1b 0 QNPN
R1  nor1q vdd 1k

*nor 2
Q3  nor2q nor2a 0 QNPN
Q4  nor2q nor2b 0 QNPN
R2  nor2q vdd 1k

*sr latch
R3  nor1q nor2a 10k
R4  nor2q nor1a 10k

* dummy loads
*R10  nor2q 0 10k     
*R11  nor1q 0 10k


.MODEL QNPN npn
+IS=1.26532e-10 BF=206.302 NF=1.5 VAF=1000
+IKF=0.0272221 ISE=2.30771e-09 NE=3.31052 BR=20.6302
+NR=2.89609 VAR=9.39809 IKR=0.272221 ISC=2.30771e-09
+NC=1.9876 RB=5.8376 IRB=50.3624 RBM=0.634251
+RE=0.0001 RC=2.65711 XTB=0.1 XTI=1
+EG=1.05 CJE=4.64214e-12 VJE=0.4 MJE=0.256227
+TF=4.19578e-10 XTF=0.906167 VTF=8.75418 ITF=0.0105823
+CJC=3.76961e-12 VJC=0.4 MJC=0.238109 XCJC=0.8
+FC=0.512134 CJS=0 VJS=0.75 MJS=0.5
+TR=6.82023e-08 PTF=0 KF=0 AF=1

.TRAN .1m 100m 

.end