VS1  VDD 0 DC 5
VS2  nor1b 0 PULSE(0 5 0 0 0 5m 20m)
VS3  nor2b 0 PULSE(0 5 10m 0 0 5m 20m)
*init sr latch
*VS4  nor1q 0 PULSE(0 5 0 0 0 1n 0)

*nor 1
Q1  nor1q nor1a 0 QNPN
Q2  nor1q nor1b 0 QNPN
R1  nor1q vdd 1k

*nor 2
Q3  nor2q nor2a 0 QNPN
Q4  nor2q nor2b 0 QNPN
R2  nor2q vdd 1k

*sr latch
R3  nor1q nor2a 10k
R4  nor2q nor1a 10k

* dummy loads
*R10  nor2q 0 10k     
*R11  nor1q 0 10k


*bc547b
.MODEL QNPN npn
+IS=7.443e-11 BF=1343.59 NF=1.42606 VAF=80.4901
+IKF=0.427163 ISE=2.4623e-10 NE=2.73946 BR=62.79
+NR=1.5 VAR=1.0092 IKR=4.27163 ISC=2.4623e-10
+NC=1.9119 RB=0.1 IRB=0.1 RBM=0.1
+RE=0.579065 RC=3.01102 XTB=0.1 XTI=2.25359
+EG=1.05 CJE=7.34106e-12 VJE=0.586136 MJE=0.33309
+TF=5.7202e-10 XTF=4.45797 VTF=26.03 ITF=0.487193
+CJC=4.04665e-12 VJC=0.95 MJC=0.343664 XCJC=0.799994
+FC=0.8 CJS=0 VJS=0.75 MJS=0.5
+TR=1e-07 PTF=0 KF=0 AF=1

.TRAN 1m 100m 

.end